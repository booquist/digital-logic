module center_light (
	input logic clk, Reset, leftLight, rightLight, leftButton, rightButton,
	output logic light
);

	logic PS, NS;
	
	parameter off = 1'b0, on = 1'b1;

	// while
	always_comb begin
		case(PS)
			off:	if (leftLight & rightButton) NS = on;           
					else if (rightLight & leftButton) NS = on;
					else NS = off;
			on:	if (rightButton | leftButton) NS = off;
					else NS = on;
			default: NS = 1'bx;	
		endcase
	end

	// reset
	always @(posedge clk)
		if (Reset)
			PS <= on; // reset should turn the center light on
		else
			PS <= NS;
			
	assign light = PS;

endmodule

module center_light_testbench();
	logic clk, Reset, leftLight, rightLight, leftButton, rightButton;
	logic light;
	
	center_light test (clk, Reset, leftLight, rightLight, leftButton, rightButton, light);
	
	// Set up a simulated clock.
	parameter CLOCK_PERIOD = 100;
	
	initial begin
		clk <= 0;
		forever #(CLOCK_PERIOD/2) clk <= ~clk; // Forever toggle the clock
	end
  
	// Set up the inputs to the design. Each line is a clock cycle.
	initial begin
		Reset <= 1;
		rightLight <= 0;
		leftLight <=0;
		leftButton <=0;
		rightButton <= 0;
		@(posedge clk);
		@(posedge clk); // Always reset FSMs at start
		Reset <= 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		leftButton <= 1;
		@(posedge clk);
		leftButton <= 0;
		@(posedge clk);
		@(posedge clk);
		leftButton <= 1;
		@(posedge clk);
		Reset <= 1;
		leftButton <= 0;
		@(posedge clk);
		Reset <= 0;
		@(posedge clk);
		rightButton <= 1;
		@(posedge clk);
		@(posedge clk);
		rightButton <= 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		Reset <= 1;
		@(posedge clk);
		leftButton <= 1;
		@(posedge clk);
		rightButton <= 1;
		$stop; // End the simulation.
	end
endmodule
	
	
	